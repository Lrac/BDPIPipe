package BDPIExample;

import BDPIPipe::*;

import "BDPI" function ActionValue#(StreamHandle) bsv_makeAdd_18b_4b;

endpackage
