package BDPIMersenneTwister;

import BDPIPipe::*;

import "BDPI" bsv_makeMersenneTwister19937 = function ActionValue#(StreamHandle) bsv_makeMersenneTwister19937;

endpackage
